`include "config.svh"

module round_robin_arbiter_with_2_requests
(
  input        clk,
  input        rst,
  input  [1:0] requests,
  output [1:0] grants
);

  // TODO: Implement the arbiter

endmodule
