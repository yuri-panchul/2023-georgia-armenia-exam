// TODO: Implement the module based on 
//
// ../03_pipelines/04_pow_5_pipelined_without_flow_control/tb.sv
// with additional flow control using signals up_rdy and down_rdy.
